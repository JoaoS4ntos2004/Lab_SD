LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY REG_BIDIRECIONAL_4B IS
  PORT(
    CLOCK    : IN  STD_LOGIC;
    RESET      : IN  STD_LOGIC;
    LOAD   : IN  STD_LOGIC;
    DADOS      : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
    DIRECAO    : IN  STD_LOGIC;
    DADO_ESQ   : IN  STD_LOGIC;
    DADO_DIR   : IN  STD_LOGIC;
    SAIDAS     : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
  );
END REG_BIDIRECIONAL_4B;

ARCHITECTURE REG_BIDIRECIONAL_4B_ARCH OF REG_BIDIRECIONAL_4B IS
  SIGNAL REGISTRO : STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
  SAIDAS <= REGISTRO;

  PROCESS(CLOCK)
  BEGIN
    IF RISING_EDGE(CLOCK) THEN
      IF RESET = '1' THEN
        REGISTRO <= (OTHERS => '0');
      ELSIF LOAD = '1' THEN
        REGISTRO <= DADOS;
      ELSIF DIRECAO = '0' THEN
        REGISTRO <= REGISTRO(2 DOWNTO 0) & DADO_ESQ;
      ELSIF DIRECAO = '1' THEN
        REGISTRO <= DADO_DIR & REGISTRO(3 DOWNTO 1);
      ELSE
        REGISTRO <= REGISTRO;
      END IF;
    END IF;
  END PROCESS;
END REG_BIDIRECIONAL_4B_ARCH;
