LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MEUCIRCUITO IS
PORT (A, B, Cin: IN STD_LOGIC;
S, Cout: OUT STD_LOGIC);
END MEUCIRCUITO;

ARCHITECTURE MEUCIRCUITO_ARCH OF MEUCIRCUITO IS
BEGIN
S <= (A XOR B) XOR Cin;
Cout <= (A AND B) OR (A AND Cin) OR (B AND Cin);
END MEUCIRCUITO_ARCH;
