LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY FLIPFLOP_JK IS
  PORT(
    PRESET   : IN  STD_LOGIC;
    CLEAR   : IN  STD_LOGIC;
    CLOCK  : IN  STD_LOGIC;
    J  : IN  STD_LOGIC;
    K : IN  STD_LOGIC;
    SAIDA    : OUT STD_LOGIC  );
END FLIPFLOP_JK;
ARCHITECTURE FLIPFLOP_JK_ARCH OF FLIPFLOP_JK IS
  SIGNAL REG : STD_LOGIC := '0';
BEGIN
   SAIDA <= REG;
 PROCESS(PRESET, CLEAR, CLOCK)
  BEGIN
    IF PRESET = '1' THEN
      REG <= '1';
    ELSIF CLEAR = '1' THEN
      REG <= '0';
    ELSIF RISING_EDGE(CLOCK) THEN
      IF J = '0' AND K = '0' THEN
        REG <= REG;
      ELSIF J = '0' AND K = '1' THEN
        REG <= '0';
      ELSIF J = '1' AND K = '0' THEN
	REG <= '1';
      ELSIF J = '1' AND K = '1' THEN
        REG <= NOT REG;
      END IF;
    END IF;
  END PROCESS;
END FLIPFLOP_JK_ARCH;
