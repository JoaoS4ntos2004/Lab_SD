LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MEUCIRCUITO2 IS
PORT (S: IN STD_LOGIC_VECTOR(0 TO 1);
D:IN STD_LOGIC_VECTOR(0 TO 3);
Y: OUT STD_LOGIC);
END MEUCIRCUITO2;

ARCHITECTURE MEUCIRCUITO2_ARCH2 OF MEUCIRCUITO2 IS
BEGIN
Y <= (D(0) AND (NOT(S(1))) AND (NOT(S(0)))) OR (D(1) AND (NOT(S(1))) 
AND S(0)) OR (D(2) AND S(1) AND (NOT(S(0)))) OR (D(3) AND S(1) AND S(0));
END MEUCIRCUITO2_ARCH2;
