LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;  
  
ENTITY SOMADOR4BIT_ARITH IS
  PORT (
    A : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
    B : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
    S : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
  );
END ENTITY;

ARCHITECTURE SOMADOR4BIT_ARITH_ARCH OF SOMADOR4BIT_ARITH IS
BEGIN
  S <= conv_std_logic_vector(
         unsigned('0' & A) + unsigned('0' & B),  
         5                                       
       );
END ARCHITECTURE SOMADOR4BIT_ARITH_ARCH;
